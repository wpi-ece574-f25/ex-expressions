module ex4(output logic [3:0] q, input logic [3:0] a, b);
    assign q = a % b;
endmodule
