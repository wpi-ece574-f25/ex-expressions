module ex2(output logic [3:0] q, input logic [1:0] a, b, c);
    assign q = a + b * c;
endmodule
