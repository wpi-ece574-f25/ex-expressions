module ex3(output logic [3:0] q, input logic [1:0] a, b);
    assign q = a + b * 2;
endmodule
